/* template_tb.v
*
* Module: module_name testbench
*
* Authors:
* author1
* author2
* author3...
*
* Description:
* This file is a template for a Verilog module testbench. The top block
* comment is strongly recommended. The rest is an example of
* organized and readble Verilog code. You may use this style if
* you wish. Regardless, make sure your code is organized and 
* neat.
*
* Revision History:
* _Rev #_	_Author(s)_	_Date_		_Changes_
* 1.00		All		mm/dd/yyyy	Module Created.
*
*/

module test ();

///////////////////////////////////////////
// Wire and Register Instantiations
//
reg [7:0] 
	8bit_reg;
reg
	reg0,
	reg1,
	reg2;
wire [7:0] 
	8bit_bus;
wire
	wire0,
	wire1,
	wire2;


template top(
	.sig1(tb_sig1),
	.sig2(tb_sig2),
	.sig3(tb_sig3)
);



endmodule // test
