/* template.v
*
* Module: module_name
*
* Authors:
* author1
* author2
* author3...
*
* Description:
* This file is a template for a Verilog module. The top block
* comment is strongly recommended. The rest is an example of
* organized and readble Verilog code. You may use this style if
* you wish. Regardless, make sure your code is organized and 
* neat.
*
* Revision History:
* _Rev #_	_Author(s)_	_Date_		_Changes_
* 1.00		All		mm/dd/yyyy	Module Created.
*
*/

// Module Declaration
module TEMPLATE (
	sig1,
	sig2,
	sig3
);

///////////////////////////////////////////
// Inputs 
//
input
	sig1,		// This is signal one
	sig2;		// This is signal two

///////////////////////////////////////////
// Outputs 
//
output
	sig3;		// This is signal three

///////////////////////////////////////////
// Wire and Register Instantiations
//
reg [7:0] 
	8bit_reg;
reg
	reg0,
	reg1,
	reg2;
wire [7:0] 
	8bit_bus;
wire
	wire0,
	wire1,
	wire2;

///////////////////////////////////////////
// YOUR LOGIC ( Use this header, as seen above )
//






endmodule // end of TEMPLATE
